PACKAGE MyPackage IS

	COMPONENT ADDER
		PORT (
			A, B, C_IN : IN BIT;
			C_OUT, S   : OUT BIT
		);
	END COMPONENT;
	
	COMPONENT FULL_ADDER
    PORT (
			VA, VB : IN  BIT_VECTOR (3 DOWNTO 0);
			VS     : OUT BIT_VECTOR (3 DOWNTO 0);
			FC_OUT : OUT BIT
		);
END COMPONENT;
   
END MyPackage;

PACKAGE BODY MyPackage IS
	CONSTANT CONSTANTE_GLOBAL: INTEGER := 200;
END MyPackage;